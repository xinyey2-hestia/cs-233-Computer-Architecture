module pipelined_machine(clk, reset);
    input        clk, reset;

    wire [31:0]  PC;
    wire [31:2]  next_PC, PC_plus4, PC_target,oldnext_PC;
    wire [31:0]  inst;

    wire [31:0]  imm = {{ 16{inst_MW[15]} }, inst_MW[15:0] };  // sign-extended immediate
    wire [4:0]   rs = inst_MW[25:21];
    wire [4:0]   rt = inst_MW[20:16];
    wire [4:0]   rd = inst_MW[15:11];
    wire [5:0]   opcode = inst_MW[31:26];
    wire [5:0]   funct = inst_MW[5:0];

    wire [4:0]   wr_regnum;
    wire [2:0]   oldALUOp,ALUOp;

    wire         RegWrite, BEQ, ALUSrc, MemRead, MemWrite, MemToReg, RegDst;
    wire         PCSrc, zero;
    wire [31:0]  rd1_data, rd2_data, B_data, alu_out_data, load_data, wr_data;

	wire  oldRegWrite, oldBEQ, oldALUSrc, oldMemRead, oldMemWrite, oldMemToReg, oldRegDst;


    // DO NOT comment out or rename this module
    // or the test bench will break
    register #(30, 30'h100000) PC_reg(PC[31:2], next_PC[31:2], clk, /* enable */~stall, reset);

    assign PC[1:0] = 2'b0;  // bottom bits hard coded to 00
    adder30 next_PC_adder(PC_plus4, PC[31:2], 30'h1);
    adder30 target_PC_adder(PC_target, PC_plus4_MW, imm[29:0]);
    mux2v #(30) branch_mux(next_PC, PC_plus4, PC_target, PCSrc);
	
    assign PCSrc = BEQ & zero;

    // DO NOT comment out or rename this module
    // or the test bench will break
    instruction_memory imem(inst, PC[31:2]);

    mips_decode decode(ALUOp, RegWrite, BEQ, ALUSrc, MemRead, MemWrite, MemToReg, RegDst,
                      opcode, funct);

    // DO NOT comment out or rename this module
    // or the test bench will break
    regfile rf (oldrd1_data, oldrd2_data,
               rs, rt, wr_regnum_MW, wr_data,
               RegWrite_MW, clk, reset);


    mux2v #(32) imm_mux(B_data, rd2_data, imm, ALUSrc);
    alu32 alu(alu_out_data, zero, ALUOp, rd1_data, B_data);

    // DO NOT comment out or rename this module
    // or the test bench will break
    data_mem data_memory(load_data, alu_out_data_MW, rd2_data_MW, MemRead_MW, MemWrite_MW, clk, reset);

    mux2v #(32) wb_mux(wr_data, alu_out_data_MW, load_data, MemToReg_MW);
    mux2v #(5) rd_mux(wr_regnum, rt, rd, RegDst);

    wire [29:0] PC_plus4_MW;
    wire [31:0] inst_MW,alu_out_data_MW,rd2_data_MW,oldrd1_data, oldrd2_data;
    wire MemRead_MW,MemWrite_MW,MemToReg_MW,RegWrite_MW;
    wire [4:0]  wr_regnum_MW;



    register #(30,30'h100000) Piplinepc (PC_plus4_MW,PC_plus4,clk,~stall,flush);
    register #(32) PiplineInstr(inst_MW,inst,clk,~stall,flush);

    register #(32) PipALUout(alu_out_data_MW,alu_out_data,clk,~stall,stall);
    register #(32) PiplineW_D(rd2_data_MW, rd2_data,clk, ~stall, stall);

    register #(1)  Piplinecontrol(MemRead_MW,MemRead,clk,~stall,stall);
  	register #(1)  Piplinecontro(MemWrite_MW,MemWrite,clk,~stall,stall);
  	register #(1)  Piplinecontr(MemToReg_MW,MemToReg,clk,~stall,stall);
	register #(1)  Piplcontr(RegWrite_MW,RegWrite,clk,~stall,stall);
  	register #(5)  Piplineconl(wr_regnum_MW,wr_regnum,clk,~stall,stall);
	
	mux2v #(32) FA(rd1_data,oldrd1_data,alu_out_data_MW,ForwardA);
	mux2v #(32) Fb(rd2_data,oldrd2_data,alu_out_data_MW,ForwardB);
	
	
	assign ForwardA = (wr_regnum_MW == rs) && RegWrite_MW&&(wr_regnum_MW!=0);
	assign ForwardB = (wr_regnum_MW == rt) && RegWrite_MW&&(wr_regnum_MW!=0);

	wire stall;

	
	assign stall = MemRead_MW && ((wr_regnum_MW == rt && RegDst) || (wr_regnum_MW == rs)) && rs != 0;
	wire flush = PCSrc || reset;
	
	


endmodule // pipelined_machine
